*ana

V1 vdd 0 3.3
V2 vin 0 1
R1 vdd vout 1000
G1 vout 0 vin 0 1
C1 vout vin 0.00000001 0
C2 vout 0 0.000001 0

.end
