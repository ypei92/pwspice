*diode

Is 0 1 1
R1 1 0 1
D1 1 0 40
D2 2 0 40
R2 1 2 1
C1 2 0 1

.end
