*Tran

V1 1 0 1
R1 2 1 1
L1 2 1 1 0
C1 2 0 1 0

.end
