*realAnalog


V1 vdd 0 3.3

V2 vin 0 1.5

M1 vout vin 0 nch 1 1

M2 vout vin vdd pch 2 1


C1 vout vin 0.00000001 0

C2 vout 0 0.000001 0



.end
