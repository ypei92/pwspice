*DC

V1 vdd 0 3.3
V2 vin 0 1
M1 vout vin 0 nch 1 1
M2 vout vin vdd pch 2 1

.end
