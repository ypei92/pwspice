*zhengliu

V1 0 xx 10
V2 1 xx 20
R1 2 0 1
D1 1 2 40

.end
