*cc
I1 1 0 1
V1 1 0 0
H1 2 0 V1 99
R1 2 0 1

.end
