*control

R1 1 0 1
Gs2 1 0 3 0 2
R3 1 2 3
R4 2 0 4
Is5 0 2 5
Vs6 3 2 6
Es7 4 0 3 0 7
R8 3 4 8

.end
